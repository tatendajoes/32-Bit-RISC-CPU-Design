`timescale 1ns/1ps

module cpu_tb;
    // Testbench for the entire CPU
    // ... Add your testbench code here ...
endmodule
