`timescale 1ns/1ps

module instruction_memory;
    // TODO: Define ports and implement instruction memory
endmodule
