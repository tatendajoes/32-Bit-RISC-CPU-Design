`timescale 1ns/1ps

module control_unit;
    // TODO: Define ports and implement control logic
endmodule
