`timescale 1ns/1ps

module design;
    // Top-level CPU design instantiating submodules
    // TODO: Connect instruction_memory, register_file, alu, control_unit, data_memory, pc
endmodule
