`timescale 1ns/1ps

module control_unit_tb;
    // Testbench for control_unit
    // ... Add your testbench code here ...
endmodule
