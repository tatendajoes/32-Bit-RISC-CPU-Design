`timescale 1ns/1ps

module instruction_memory_tb;
    // Testbench for instruction_memory
    // ... Add your testbench code here ...
endmodule
